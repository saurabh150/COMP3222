library verilog;
use verilog.vl_types.all;
entity L2P21_vlg_vec_tst is
end L2P21_vlg_vec_tst;
