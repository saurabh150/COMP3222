LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY L1P1 IS
	PORT (SW		:IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
			Ledr	:OUT	STD_LOGIC_VECTOR(9 DOWNTO 0));
END L1P1;

ARCHITECTURE Behavior OF L1P1 IS
BEGIN
	LEDR <= SW;
END Behavior;