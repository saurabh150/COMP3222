library verilog;
use verilog.vl_types.all;
entity L4P1_vlg_vec_tst is
end L4P1_vlg_vec_tst;
