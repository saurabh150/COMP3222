LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY L1P2 IS 
PORT (SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
      LEDG : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END L1P2;

ARCHITECTURE Behavior OF L1P2 IS
SIGNAL	X: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	Y:	STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	S:	STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	M: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	X<=SW(3 DOWNTO 0);
	Y<=SW(7 DOWNTO 4);
	S(0)<=SW(9);
	S(1)<=SW(9);
	S(2)<=SW(9);
	S(3)<=SW(9);
	M<=(NOT S AND X) OR (S AND Y);
	LEDG<=M;
	
END Behavior;
